module Test();
endmodule
